`timescale 1ns / 1ps

// charmap.vpp 
// module to map the a character given on the input, together with a pixel offset, into a binary pixel value. 
// done by a lookup table ( a ROM). 

// ports: 

// CLK_108MHz - global clock

// reset - global, async, reset

// hctr_in - horixontal pixel value. 3 bits. 

// vctr_in - vertical pixel value. 3 bits. 

// character_in - what character it is. 8 bits. 

// color_in - used in the next stage to give the colored output, so register. 8 bits. 

// hsync_in - hsync, needs registred

// vsync_in - vsync, needs registred

// de_in - de, needs registred. 

// pixel_out - the value of the pixel. 

// color_out - color output for the next stage

// hsync_out - registred hsync value

// vsync_out - registred vsync value

// de_out - registred de value


module charmap(

input CLK_108MHz,
input reset,
input [2:0] hctr_in,
input [2:0] vctr_in,
input [7:0] character_in,
input [7:0] color_in,
input hsync_in,
input vsync_in,
input de_in,
output reg pixel_out,
output reg [7:0] color_out,
output reg hsync_out,
output reg vsync_out,
output reg de_out
);

reg [8191:0] charmap;

initial begin

charmap [7:0]  = 8'b00000000;
charmap [15:8]  = 8'b00000000;
charmap [23:16]  = 8'b00000000;
charmap [31:24]  = 8'b00000000;
charmap [39:32]  = 8'b00000000;
charmap [47:40]  = 8'b00000000;
charmap [55:48]  = 8'b00000000;
charmap [63:56]  = 8'b00000000;
charmap [71:64]  = 8'b00011100;
charmap [79:72]  = 8'b00100010;
charmap [87:80]  = 8'b00100010;
charmap [95:88]  = 8'b00101010;
charmap [103:96]  = 8'b00100010;
charmap [111:104]  = 8'b00100010;
charmap [119:112]  = 8'b00011100;
charmap [127:120]  = 8'b00000000;
charmap [135:128]  = 8'b00000000;
charmap [143:136]  = 8'b00000000;
charmap [151:144]  = 8'b00000000;
charmap [159:152]  = 8'b00000000;
charmap [167:160]  = 8'b00000000;
charmap [175:168]  = 8'b00000000;
charmap [183:176]  = 8'b00000000;
charmap [191:184]  = 8'b00000000;
charmap [199:192]  = 8'b00001000;
charmap [207:200]  = 8'b00001100;
charmap [215:208]  = 8'b00001000;
charmap [223:216]  = 8'b00001000;
charmap [231:224]  = 8'b00001000;
charmap [239:232]  = 8'b00001000;
charmap [247:240]  = 8'b00011100;
charmap [255:248]  = 8'b00000000;
charmap [263:256]  = 8'b00000000;
charmap [271:264]  = 8'b00000000;
charmap [279:272]  = 8'b00000000;
charmap [287:280]  = 8'b00000000;
charmap [295:288]  = 8'b00000000;
charmap [303:296]  = 8'b00000000;
charmap [311:304]  = 8'b00000000;
charmap [319:312]  = 8'b00000000;
charmap [327:320]  = 8'b00011100;
charmap [335:328]  = 8'b00100010;
charmap [343:336]  = 8'b00100000;
charmap [351:344]  = 8'b00010000;
charmap [359:352]  = 8'b00001000;
charmap [367:360]  = 8'b00000100;
charmap [375:368]  = 8'b00111110;
charmap [383:376]  = 8'b00000000;
charmap [391:384]  = 8'b00000000;
charmap [399:392]  = 8'b00000000;
charmap [407:400]  = 8'b00000000;
charmap [415:408]  = 8'b00000000;
charmap [423:416]  = 8'b00000000;
charmap [431:424]  = 8'b00000000;
charmap [439:432]  = 8'b00000000;
charmap [447:440]  = 8'b00000000;
charmap [455:448]  = 8'b00011100;
charmap [463:456]  = 8'b00100010;
charmap [471:464]  = 8'b00100000;
charmap [479:472]  = 8'b00011000;
charmap [487:480]  = 8'b00100000;
charmap [495:488]  = 8'b00100010;
charmap [503:496]  = 8'b00011100;
charmap [511:504]  = 8'b00000000;
charmap [519:512]  = 8'b00000000;
charmap [527:520]  = 8'b00000000;
charmap [535:528]  = 8'b00000000;
charmap [543:536]  = 8'b00000000;
charmap [551:544]  = 8'b00000000;
charmap [559:552]  = 8'b00000000;
charmap [567:560]  = 8'b00000000;
charmap [575:568]  = 8'b00000000;
charmap [583:576]  = 8'b00001000;
charmap [591:584]  = 8'b00010000;
charmap [599:592]  = 8'b00100000;
charmap [607:600]  = 8'b01111110;
charmap [615:608]  = 8'b00100000;
charmap [623:616]  = 8'b00010000;
charmap [631:624]  = 8'b00001000;
charmap [639:632]  = 8'b00000000;
charmap [647:640]  = 8'b00000000;
charmap [655:648]  = 8'b00000000;
charmap [663:656]  = 8'b00000000;
charmap [671:664]  = 8'b00000000;
charmap [679:672]  = 8'b00000000;
charmap [687:680]  = 8'b00000000;
charmap [695:688]  = 8'b00000000;
charmap [703:696]  = 8'b00000000;
charmap [711:704]  = 8'b00111110;
charmap [719:712]  = 8'b00000010;
charmap [727:720]  = 8'b00000010;
charmap [735:728]  = 8'b00011110;
charmap [743:736]  = 8'b00100000;
charmap [751:744]  = 8'b00100010;
charmap [759:752]  = 8'b00011100;
charmap [767:760]  = 8'b00000000;
charmap [775:768]  = 8'b00000000;
charmap [783:776]  = 8'b00000000;
charmap [791:784]  = 8'b00000000;
charmap [799:792]  = 8'b00000000;
charmap [807:800]  = 8'b00000000;
charmap [815:808]  = 8'b00000000;
charmap [823:816]  = 8'b00000000;
charmap [831:824]  = 8'b00000000;
charmap [839:832]  = 8'b00000000;
charmap [847:840]  = 8'b00000000;
charmap [855:848]  = 8'b00000000;
charmap [863:856]  = 8'b00000000;
charmap [871:864]  = 8'b00000000;
charmap [879:872]  = 8'b00000000;
charmap [887:880]  = 8'b00000000;
charmap [895:888]  = 8'b00000000;
charmap [903:896]  = 8'b00000000;
charmap [911:904]  = 8'b00000000;
charmap [919:912]  = 8'b00000000;
charmap [927:920]  = 8'b00000000;
charmap [935:928]  = 8'b00000000;
charmap [943:936]  = 8'b00000000;
charmap [951:944]  = 8'b00000000;
charmap [959:952]  = 8'b00000000;
charmap [967:960]  = 8'b00111110;
charmap [975:968]  = 8'b00100000;
charmap [983:976]  = 8'b00010000;
charmap [991:984]  = 8'b00001000;
charmap [999:992]  = 8'b00000100;
charmap [1007:1000]  = 8'b00000100;
charmap [1015:1008]  = 8'b00000100;
charmap [1023:1016]  = 8'b00000000;
charmap [1031:1024]  = 8'b00000000;
charmap [1039:1032]  = 8'b00000000;
charmap [1047:1040]  = 8'b00000000;
charmap [1055:1048]  = 8'b00000000;
charmap [1063:1056]  = 8'b00000000;
charmap [1071:1064]  = 8'b00000000;
charmap [1079:1072]  = 8'b00000000;
charmap [1087:1080]  = 8'b00000000;
charmap [1095:1088]  = 8'b00011100;
charmap [1103:1096]  = 8'b00100010;
charmap [1111:1104]  = 8'b00100010;
charmap [1119:1112]  = 8'b00011100;
charmap [1127:1120]  = 8'b00100010;
charmap [1135:1128]  = 8'b00100010;
charmap [1143:1136]  = 8'b00011100;
charmap [1151:1144]  = 8'b00000000;
charmap [1159:1152]  = 8'b00000000;
charmap [1167:1160]  = 8'b00000000;
charmap [1175:1168]  = 8'b00000000;
charmap [1183:1176]  = 8'b00000000;
charmap [1191:1184]  = 8'b00000000;
charmap [1199:1192]  = 8'b00000000;
charmap [1207:1200]  = 8'b00000000;
charmap [1215:1208]  = 8'b00000000;
charmap [1223:1216]  = 8'b00011100;
charmap [1231:1224]  = 8'b00100010;
charmap [1239:1232]  = 8'b00100010;
charmap [1247:1240]  = 8'b00111100;
charmap [1255:1248]  = 8'b00100000;
charmap [1263:1256]  = 8'b00100010;
charmap [1271:1264]  = 8'b00011100;
charmap [1279:1272]  = 8'b00000000;
charmap [1287:1280]  = 8'b00000000;
charmap [1295:1288]  = 8'b00000000;
charmap [1303:1296]  = 8'b00000000;
charmap [1311:1304]  = 8'b00000000;
charmap [1319:1312]  = 8'b00000000;
charmap [1327:1320]  = 8'b00000000;
charmap [1335:1328]  = 8'b00000000;
charmap [1343:1336]  = 8'b00000000;
charmap [1351:1344]  = 8'b00011100;
charmap [1359:1352]  = 8'b00100010;
charmap [1367:1360]  = 8'b00100010;
charmap [1375:1368]  = 8'b00111110;
charmap [1383:1376]  = 8'b00100010;
charmap [1391:1384]  = 8'b00100010;
charmap [1399:1392]  = 8'b00100010;
charmap [1407:1400]  = 8'b00000000;
charmap [1415:1408]  = 8'b00000000;
charmap [1423:1416]  = 8'b00000000;
charmap [1431:1424]  = 8'b00000000;
charmap [1439:1432]  = 8'b00000000;
charmap [1447:1440]  = 8'b00000000;
charmap [1455:1448]  = 8'b00000000;
charmap [1463:1456]  = 8'b00000000;
charmap [1471:1464]  = 8'b00000000;
charmap [1479:1472]  = 8'b00011110;
charmap [1487:1480]  = 8'b00100010;
charmap [1495:1488]  = 8'b00100010;
charmap [1503:1496]  = 8'b00011110;
charmap [1511:1504]  = 8'b00100010;
charmap [1519:1512]  = 8'b00100010;
charmap [1527:1520]  = 8'b00011110;
charmap [1535:1528]  = 8'b00000000;
charmap [1543:1536]  = 8'b00000000;
charmap [1551:1544]  = 8'b00000000;
charmap [1559:1552]  = 8'b00000000;
charmap [1567:1560]  = 8'b00000000;
charmap [1575:1568]  = 8'b00000000;
charmap [1583:1576]  = 8'b00000000;
charmap [1591:1584]  = 8'b00000000;
charmap [1599:1592]  = 8'b00000000;
charmap [1607:1600]  = 8'b00011100;
charmap [1615:1608]  = 8'b00100010;
charmap [1623:1616]  = 8'b00000010;
charmap [1631:1624]  = 8'b00000010;
charmap [1639:1632]  = 8'b00000010;
charmap [1647:1640]  = 8'b00100010;
charmap [1655:1648]  = 8'b00011100;
charmap [1663:1656]  = 8'b00000000;
charmap [1671:1664]  = 8'b00000000;
charmap [1679:1672]  = 8'b00000000;
charmap [1687:1680]  = 8'b00000000;
charmap [1695:1688]  = 8'b00000000;
charmap [1703:1696]  = 8'b00000000;
charmap [1711:1704]  = 8'b00000000;
charmap [1719:1712]  = 8'b00000000;
charmap [1727:1720]  = 8'b00000000;
charmap [1735:1728]  = 8'b00011110;
charmap [1743:1736]  = 8'b00100010;
charmap [1751:1744]  = 8'b00100010;
charmap [1759:1752]  = 8'b00100010;
charmap [1767:1760]  = 8'b00100010;
charmap [1775:1768]  = 8'b00100010;
charmap [1783:1776]  = 8'b00011110;
charmap [1791:1784]  = 8'b00000000;
charmap [1799:1792]  = 8'b00000000;
charmap [1807:1800]  = 8'b00000000;
charmap [1815:1808]  = 8'b00000000;
charmap [1823:1816]  = 8'b00000000;
charmap [1831:1824]  = 8'b00000000;
charmap [1839:1832]  = 8'b00000000;
charmap [1847:1840]  = 8'b00000000;
charmap [1855:1848]  = 8'b00000000;
charmap [1863:1856]  = 8'b00111110;
charmap [1871:1864]  = 8'b00000010;
charmap [1879:1872]  = 8'b00000010;
charmap [1887:1880]  = 8'b00011110;
charmap [1895:1888]  = 8'b00000010;
charmap [1903:1896]  = 8'b00000010;
charmap [1911:1904]  = 8'b00111110;
charmap [1919:1912]  = 8'b00000000;
charmap [1927:1920]  = 8'b00000000;
charmap [1935:1928]  = 8'b00000000;
charmap [1943:1936]  = 8'b00000000;
charmap [1951:1944]  = 8'b00000000;
charmap [1959:1952]  = 8'b00000000;
charmap [1967:1960]  = 8'b00000000;
charmap [1975:1968]  = 8'b00000000;
charmap [1983:1976]  = 8'b00000000;
charmap [1991:1984]  = 8'b00111110;
charmap [1999:1992]  = 8'b00000010;
charmap [2007:2000]  = 8'b00000010;
charmap [2015:2008]  = 8'b00111110;
charmap [2023:2016]  = 8'b00000010;
charmap [2031:2024]  = 8'b00000010;
charmap [2039:2032]  = 8'b00000010;
charmap [2047:2040]  = 8'b00000000;
charmap [2055:2048]  = 8'b00000000;
charmap [2063:2056]  = 8'b00000000;
charmap [2071:2064]  = 8'b00000000;
charmap [2079:2072]  = 8'b00000000;
charmap [2087:2080]  = 8'b00000000;
charmap [2095:2088]  = 8'b00000000;
charmap [2103:2096]  = 8'b00000000;
charmap [2111:2104]  = 8'b00000000;
charmap [2119:2112]  = 8'b00010000;
charmap [2127:2120]  = 8'b00010000;
charmap [2135:2128]  = 8'b00010000;
charmap [2143:2136]  = 8'b00010000;
charmap [2151:2144]  = 8'b00010000;
charmap [2159:2152]  = 8'b00000000;
charmap [2167:2160]  = 8'b00010000;
charmap [2175:2168]  = 8'b00000000;
charmap [2183:2176]  = 8'b00101000;
charmap [2191:2184]  = 8'b00101000;
charmap [2199:2192]  = 8'b00000000;
charmap [2207:2200]  = 8'b00000000;
charmap [2215:2208]  = 8'b00000000;
charmap [2223:2216]  = 8'b00000000;
charmap [2231:2224]  = 8'b00000000;
charmap [2239:2232]  = 8'b00000000;
charmap [2247:2240]  = 8'b00101000;
charmap [2255:2248]  = 8'b00101000;
charmap [2263:2256]  = 8'b11111110;
charmap [2271:2264]  = 8'b00101000;
charmap [2279:2272]  = 8'b11111110;
charmap [2287:2280]  = 8'b00101000;
charmap [2295:2288]  = 8'b00101000;
charmap [2303:2296]  = 8'b00000000;
charmap [2311:2304]  = 8'b00010000;
charmap [2319:2312]  = 8'b01111000;
charmap [2327:2320]  = 8'b00010100;
charmap [2335:2328]  = 8'b00111000;
charmap [2343:2336]  = 8'b01010000;
charmap [2351:2344]  = 8'b00111100;
charmap [2359:2352]  = 8'b00010000;
charmap [2367:2360]  = 8'b00000000;
charmap [2375:2368]  = 8'b00000000;
charmap [2383:2376]  = 8'b01001100;
charmap [2391:2384]  = 8'b00101100;
charmap [2399:2392]  = 8'b00010000;
charmap [2407:2400]  = 8'b01101000;
charmap [2415:2408]  = 8'b01100100;
charmap [2423:2416]  = 8'b00000000;
charmap [2431:2424]  = 8'b00000000;
charmap [2439:2432]  = 8'b00011000;
charmap [2447:2440]  = 8'b00010100;
charmap [2455:2448]  = 8'b00001000;
charmap [2463:2456]  = 8'b00010100;
charmap [2471:2464]  = 8'b01100010;
charmap [2479:2472]  = 8'b00100010;
charmap [2487:2480]  = 8'b01011100;
charmap [2495:2488]  = 8'b00000000;
charmap [2503:2496]  = 8'b00010000;
charmap [2511:2504]  = 8'b00010000;
charmap [2519:2512]  = 8'b00000000;
charmap [2527:2520]  = 8'b00000000;
charmap [2535:2528]  = 8'b00000000;
charmap [2543:2536]  = 8'b00000000;
charmap [2551:2544]  = 8'b00000000;
charmap [2559:2552]  = 8'b00000000;
charmap [2567:2560]  = 8'b00100000;
charmap [2575:2568]  = 8'b00010000;
charmap [2583:2576]  = 8'b00001000;
charmap [2591:2584]  = 8'b00001000;
charmap [2599:2592]  = 8'b00001000;
charmap [2607:2600]  = 8'b00010000;
charmap [2615:2608]  = 8'b00100000;
charmap [2623:2616]  = 8'b00000000;
charmap [2631:2624]  = 8'b00001000;
charmap [2639:2632]  = 8'b00010000;
charmap [2647:2640]  = 8'b00100000;
charmap [2655:2648]  = 8'b00100000;
charmap [2663:2656]  = 8'b00100000;
charmap [2671:2664]  = 8'b00010000;
charmap [2679:2672]  = 8'b00001000;
charmap [2687:2680]  = 8'b00000000;
charmap [2695:2688]  = 8'b00010000;
charmap [2703:2696]  = 8'b10010010;
charmap [2711:2704]  = 8'b01010100;
charmap [2719:2712]  = 8'b00111000;
charmap [2727:2720]  = 8'b01010100;
charmap [2735:2728]  = 8'b10010010;
charmap [2743:2736]  = 8'b00010000;
charmap [2751:2744]  = 8'b00000000;
charmap [2759:2752]  = 8'b00010000;
charmap [2767:2760]  = 8'b00010000;
charmap [2775:2768]  = 8'b00010000;
charmap [2783:2776]  = 8'b11111110;
charmap [2791:2784]  = 8'b00010000;
charmap [2799:2792]  = 8'b00010000;
charmap [2807:2800]  = 8'b00010000;
charmap [2815:2808]  = 8'b00000000;
charmap [2823:2816]  = 8'b00000000;
charmap [2831:2824]  = 8'b00000000;
charmap [2839:2832]  = 8'b00000000;
charmap [2847:2840]  = 8'b00000000;
charmap [2855:2848]  = 8'b00110000;
charmap [2863:2856]  = 8'b00110000;
charmap [2871:2864]  = 8'b00100000;
charmap [2879:2872]  = 8'b00010000;
charmap [2887:2880]  = 8'b00000000;
charmap [2895:2888]  = 8'b00000000;
charmap [2903:2896]  = 8'b00000000;
charmap [2911:2904]  = 8'b11111110;
charmap [2919:2912]  = 8'b00000000;
charmap [2927:2920]  = 8'b00000000;
charmap [2935:2928]  = 8'b00000000;
charmap [2943:2936]  = 8'b00000000;
charmap [2951:2944]  = 8'b00000000;
charmap [2959:2952]  = 8'b00000000;
charmap [2967:2960]  = 8'b00000000;
charmap [2975:2968]  = 8'b00000000;
charmap [2983:2976]  = 8'b00000000;
charmap [2991:2984]  = 8'b00110000;
charmap [2999:2992]  = 8'b00110000;
charmap [3007:3000]  = 8'b00000000;
charmap [3015:3008]  = 8'b10000000;
charmap [3023:3016]  = 8'b01000000;
charmap [3031:3024]  = 8'b00100000;
charmap [3039:3032]  = 8'b00010000;
charmap [3047:3040]  = 8'b00001000;
charmap [3055:3048]  = 8'b00000100;
charmap [3063:3056]  = 8'b00000010;
charmap [3071:3064]  = 8'b00000000;
charmap [3079:3072]  = 8'b00111000;
charmap [3087:3080]  = 8'b01000100;
charmap [3095:3088]  = 8'b01000100;
charmap [3103:3096]  = 8'b01010100;
charmap [3111:3104]  = 8'b01000100;
charmap [3119:3112]  = 8'b01000100;
charmap [3127:3120]  = 8'b00111000;
charmap [3135:3128]  = 8'b00000000;
charmap [3143:3136]  = 8'b00010000;
charmap [3151:3144]  = 8'b00011000;
charmap [3159:3152]  = 8'b00010000;
charmap [3167:3160]  = 8'b00010000;
charmap [3175:3168]  = 8'b00010000;
charmap [3183:3176]  = 8'b00010000;
charmap [3191:3184]  = 8'b00111000;
charmap [3199:3192]  = 8'b00000000;
charmap [3207:3200]  = 8'b00111000;
charmap [3215:3208]  = 8'b01000100;
charmap [3223:3216]  = 8'b01000000;
charmap [3231:3224]  = 8'b00100000;
charmap [3239:3232]  = 8'b00010000;
charmap [3247:3240]  = 8'b00001000;
charmap [3255:3248]  = 8'b01111100;
charmap [3263:3256]  = 8'b00000000;
charmap [3271:3264]  = 8'b00111000;
charmap [3279:3272]  = 8'b01000100;
charmap [3287:3280]  = 8'b01000000;
charmap [3295:3288]  = 8'b00110000;
charmap [3303:3296]  = 8'b01000000;
charmap [3311:3304]  = 8'b01000100;
charmap [3319:3312]  = 8'b00111000;
charmap [3327:3320]  = 8'b00000000;
charmap [3335:3328]  = 8'b00110000;
charmap [3343:3336]  = 8'b00101000;
charmap [3351:3344]  = 8'b00100100;
charmap [3359:3352]  = 8'b01111100;
charmap [3367:3360]  = 8'b00100000;
charmap [3375:3368]  = 8'b00100000;
charmap [3383:3376]  = 8'b01110000;
charmap [3391:3384]  = 8'b00000000;
charmap [3399:3392]  = 8'b01111100;
charmap [3407:3400]  = 8'b00000100;
charmap [3415:3408]  = 8'b00000100;
charmap [3423:3416]  = 8'b00111100;
charmap [3431:3424]  = 8'b01000000;
charmap [3439:3432]  = 8'b01000100;
charmap [3447:3440]  = 8'b00111000;
charmap [3455:3448]  = 8'b00000000;
charmap [3463:3456]  = 8'b00111000;
charmap [3471:3464]  = 8'b01000100;
charmap [3479:3472]  = 8'b00000100;
charmap [3487:3480]  = 8'b00111100;
charmap [3495:3488]  = 8'b01000100;
charmap [3503:3496]  = 8'b01000100;
charmap [3511:3504]  = 8'b00111000;
charmap [3519:3512]  = 8'b00000000;
charmap [3527:3520]  = 8'b01111100;
charmap [3535:3528]  = 8'b01000000;
charmap [3543:3536]  = 8'b00100000;
charmap [3551:3544]  = 8'b00010000;
charmap [3559:3552]  = 8'b00001000;
charmap [3567:3560]  = 8'b00001000;
charmap [3575:3568]  = 8'b00001000;
charmap [3583:3576]  = 8'b00000000;
charmap [3591:3584]  = 8'b00111000;
charmap [3599:3592]  = 8'b01000100;
charmap [3607:3600]  = 8'b01000100;
charmap [3615:3608]  = 8'b00111000;
charmap [3623:3616]  = 8'b01000100;
charmap [3631:3624]  = 8'b01000100;
charmap [3639:3632]  = 8'b00111000;
charmap [3647:3640]  = 8'b00000000;
charmap [3655:3648]  = 8'b00111000;
charmap [3663:3656]  = 8'b01000100;
charmap [3671:3664]  = 8'b01000100;
charmap [3679:3672]  = 8'b01111000;
charmap [3687:3680]  = 8'b01000000;
charmap [3695:3688]  = 8'b01000100;
charmap [3703:3696]  = 8'b00111000;
charmap [3711:3704]  = 8'b00000000;
charmap [3719:3712]  = 8'b00000000;
charmap [3727:3720]  = 8'b00110000;
charmap [3735:3728]  = 8'b00110000;
charmap [3743:3736]  = 8'b00000000;
charmap [3751:3744]  = 8'b00110000;
charmap [3759:3752]  = 8'b00110000;
charmap [3767:3760]  = 8'b00000000;
charmap [3775:3768]  = 8'b00000000;
charmap [3783:3776]  = 8'b00000000;
charmap [3791:3784]  = 8'b00110000;
charmap [3799:3792]  = 8'b00110000;
charmap [3807:3800]  = 8'b00000000;
charmap [3815:3808]  = 8'b00110000;
charmap [3823:3816]  = 8'b00110000;
charmap [3831:3824]  = 8'b00100000;
charmap [3839:3832]  = 8'b00010000;
charmap [3847:3840]  = 8'b00100000;
charmap [3855:3848]  = 8'b00010000;
charmap [3863:3856]  = 8'b00001000;
charmap [3871:3864]  = 8'b00000100;
charmap [3879:3872]  = 8'b00001000;
charmap [3887:3880]  = 8'b00010000;
charmap [3895:3888]  = 8'b00100000;
charmap [3903:3896]  = 8'b00000000;
charmap [3911:3904]  = 8'b00000000;
charmap [3919:3912]  = 8'b00000000;
charmap [3927:3920]  = 8'b11111110;
charmap [3935:3928]  = 8'b00000000;
charmap [3943:3936]  = 8'b11111110;
charmap [3951:3944]  = 8'b00000000;
charmap [3959:3952]  = 8'b00000000;
charmap [3967:3960]  = 8'b00000000;
charmap [3975:3968]  = 8'b00000100;
charmap [3983:3976]  = 8'b00001000;
charmap [3991:3984]  = 8'b00010000;
charmap [3999:3992]  = 8'b00100000;
charmap [4007:4000]  = 8'b00010000;
charmap [4015:4008]  = 8'b00001000;
charmap [4023:4016]  = 8'b00000100;
charmap [4031:4024]  = 8'b00000000;
charmap [4039:4032]  = 8'b00111000;
charmap [4047:4040]  = 8'b01000100;
charmap [4055:4048]  = 8'b01000000;
charmap [4063:4056]  = 8'b00100000;
charmap [4071:4064]  = 8'b00010000;
charmap [4079:4072]  = 8'b00000000;
charmap [4087:4080]  = 8'b00010000;
charmap [4095:4088]  = 8'b00000000;
charmap [4103:4096]  = 8'b00111000;
charmap [4111:4104]  = 8'b01000100;
charmap [4119:4112]  = 8'b01110100;
charmap [4127:4120]  = 8'b01010100;
charmap [4135:4128]  = 8'b01110100;
charmap [4143:4136]  = 8'b00000100;
charmap [4151:4144]  = 8'b00111000;
charmap [4159:4152]  = 8'b00000000;
charmap [4167:4160]  = 8'b00111000;
charmap [4175:4168]  = 8'b01000100;
charmap [4183:4176]  = 8'b01000100;
charmap [4191:4184]  = 8'b01111100;
charmap [4199:4192]  = 8'b01000100;
charmap [4207:4200]  = 8'b01000100;
charmap [4215:4208]  = 8'b01000100;
charmap [4223:4216]  = 8'b00000000;
charmap [4231:4224]  = 8'b00111100;
charmap [4239:4232]  = 8'b01000100;
charmap [4247:4240]  = 8'b01000100;
charmap [4255:4248]  = 8'b00111100;
charmap [4263:4256]  = 8'b01000100;
charmap [4271:4264]  = 8'b01000100;
charmap [4279:4272]  = 8'b00111100;
charmap [4287:4280]  = 8'b00000000;
charmap [4295:4288]  = 8'b00111000;
charmap [4303:4296]  = 8'b01000100;
charmap [4311:4304]  = 8'b00000100;
charmap [4319:4312]  = 8'b00000100;
charmap [4327:4320]  = 8'b00000100;
charmap [4335:4328]  = 8'b01000100;
charmap [4343:4336]  = 8'b00111000;
charmap [4351:4344]  = 8'b00000000;
charmap [4359:4352]  = 8'b00111100;
charmap [4367:4360]  = 8'b01000100;
charmap [4375:4368]  = 8'b01000100;
charmap [4383:4376]  = 8'b01000100;
charmap [4391:4384]  = 8'b01000100;
charmap [4399:4392]  = 8'b01000100;
charmap [4407:4400]  = 8'b00111100;
charmap [4415:4408]  = 8'b00000000;
charmap [4423:4416]  = 8'b01111100;
charmap [4431:4424]  = 8'b00000100;
charmap [4439:4432]  = 8'b00000100;
charmap [4447:4440]  = 8'b00111100;
charmap [4455:4448]  = 8'b00000100;
charmap [4463:4456]  = 8'b00000100;
charmap [4471:4464]  = 8'b01111100;
charmap [4479:4472]  = 8'b00000000;
charmap [4487:4480]  = 8'b01111100;
charmap [4495:4488]  = 8'b00000100;
charmap [4503:4496]  = 8'b00000100;
charmap [4511:4504]  = 8'b01111100;
charmap [4519:4512]  = 8'b00000100;
charmap [4527:4520]  = 8'b00000100;
charmap [4535:4528]  = 8'b00000100;
charmap [4543:4536]  = 8'b00000000;
charmap [4551:4544]  = 8'b00111000;
charmap [4559:4552]  = 8'b01000100;
charmap [4567:4560]  = 8'b00000100;
charmap [4575:4568]  = 8'b01110100;
charmap [4583:4576]  = 8'b01000100;
charmap [4591:4584]  = 8'b01000100;
charmap [4599:4592]  = 8'b00111000;
charmap [4607:4600]  = 8'b00000000;
charmap [4615:4608]  = 8'b01000100;
charmap [4623:4616]  = 8'b01000100;
charmap [4631:4624]  = 8'b01000100;
charmap [4639:4632]  = 8'b01111100;
charmap [4647:4640]  = 8'b01000100;
charmap [4655:4648]  = 8'b01000100;
charmap [4663:4656]  = 8'b01000100;
charmap [4671:4664]  = 8'b00000000;
charmap [4679:4672]  = 8'b00111000;
charmap [4687:4680]  = 8'b00010000;
charmap [4695:4688]  = 8'b00010000;
charmap [4703:4696]  = 8'b00010000;
charmap [4711:4704]  = 8'b00010000;
charmap [4719:4712]  = 8'b00010000;
charmap [4727:4720]  = 8'b00111000;
charmap [4735:4728]  = 8'b00000000;
charmap [4743:4736]  = 8'b01110000;
charmap [4751:4744]  = 8'b00100000;
charmap [4759:4752]  = 8'b00100000;
charmap [4767:4760]  = 8'b00100000;
charmap [4775:4768]  = 8'b00100100;
charmap [4783:4776]  = 8'b00100100;
charmap [4791:4784]  = 8'b00011000;
charmap [4799:4792]  = 8'b00000000;
charmap [4807:4800]  = 8'b01000100;
charmap [4815:4808]  = 8'b01000100;
charmap [4823:4816]  = 8'b00100100;
charmap [4831:4824]  = 8'b00011100;
charmap [4839:4832]  = 8'b00100100;
charmap [4847:4840]  = 8'b01000100;
charmap [4855:4848]  = 8'b01000100;
charmap [4863:4856]  = 8'b00000000;
charmap [4871:4864]  = 8'b00001000;
charmap [4879:4872]  = 8'b00001000;
charmap [4887:4880]  = 8'b00001000;
charmap [4895:4888]  = 8'b00001000;
charmap [4903:4896]  = 8'b00001000;
charmap [4911:4904]  = 8'b00001000;
charmap [4919:4912]  = 8'b01111000;
charmap [4927:4920]  = 8'b00000000;
charmap [4935:4928]  = 8'b10000010;
charmap [4943:4936]  = 8'b11000110;
charmap [4951:4944]  = 8'b10101010;
charmap [4959:4952]  = 8'b10010010;
charmap [4967:4960]  = 8'b10000010;
charmap [4975:4968]  = 8'b10000010;
charmap [4983:4976]  = 8'b10000010;
charmap [4991:4984]  = 8'b00000000;
charmap [4999:4992]  = 8'b01000100;
charmap [5007:5000]  = 8'b01001100;
charmap [5015:5008]  = 8'b01010100;
charmap [5023:5016]  = 8'b01010100;
charmap [5031:5024]  = 8'b01100100;
charmap [5039:5032]  = 8'b01000100;
charmap [5047:5040]  = 8'b01000100;
charmap [5055:5048]  = 8'b00000000;
charmap [5063:5056]  = 8'b00111000;
charmap [5071:5064]  = 8'b01000100;
charmap [5079:5072]  = 8'b01000100;
charmap [5087:5080]  = 8'b01000100;
charmap [5095:5088]  = 8'b01000100;
charmap [5103:5096]  = 8'b01000100;
charmap [5111:5104]  = 8'b00111000;
charmap [5119:5112]  = 8'b00000000;
charmap [5127:5120]  = 8'b00111000;
charmap [5135:5128]  = 8'b01001000;
charmap [5143:5136]  = 8'b01001000;
charmap [5151:5144]  = 8'b00111000;
charmap [5159:5152]  = 8'b00001000;
charmap [5167:5160]  = 8'b00001000;
charmap [5175:5168]  = 8'b00001000;
charmap [5183:5176]  = 8'b00000000;
charmap [5191:5184]  = 8'b00111000;
charmap [5199:5192]  = 8'b01000100;
charmap [5207:5200]  = 8'b01000100;
charmap [5215:5208]  = 8'b01000100;
charmap [5223:5216]  = 8'b01000100;
charmap [5231:5224]  = 8'b01000100;
charmap [5239:5232]  = 8'b00111000;
charmap [5247:5240]  = 8'b01100000;
charmap [5255:5248]  = 8'b00111100;
charmap [5263:5256]  = 8'b01000100;
charmap [5271:5264]  = 8'b01000100;
charmap [5279:5272]  = 8'b00111100;
charmap [5287:5280]  = 8'b00010100;
charmap [5295:5288]  = 8'b00100100;
charmap [5303:5296]  = 8'b01000100;
charmap [5311:5304]  = 8'b00000000;
charmap [5319:5312]  = 8'b00111000;
charmap [5327:5320]  = 8'b01000100;
charmap [5335:5328]  = 8'b00000100;
charmap [5343:5336]  = 8'b00111000;
charmap [5351:5344]  = 8'b01000000;
charmap [5359:5352]  = 8'b01000100;
charmap [5367:5360]  = 8'b00111000;
charmap [5375:5368]  = 8'b00000000;
charmap [5383:5376]  = 8'b01111100;
charmap [5391:5384]  = 8'b00010000;
charmap [5399:5392]  = 8'b00010000;
charmap [5407:5400]  = 8'b00010000;
charmap [5415:5408]  = 8'b00010000;
charmap [5423:5416]  = 8'b00010000;
charmap [5431:5424]  = 8'b00010000;
charmap [5439:5432]  = 8'b00000000;
charmap [5447:5440]  = 8'b01000100;
charmap [5455:5448]  = 8'b01000100;
charmap [5463:5456]  = 8'b01000100;
charmap [5471:5464]  = 8'b01000100;
charmap [5479:5472]  = 8'b01000100;
charmap [5487:5480]  = 8'b01000100;
charmap [5495:5488]  = 8'b00111000;
charmap [5503:5496]  = 8'b00000000;
charmap [5511:5504]  = 8'b01000100;
charmap [5519:5512]  = 8'b01000100;
charmap [5527:5520]  = 8'b01000100;
charmap [5535:5528]  = 8'b00101000;
charmap [5543:5536]  = 8'b00101000;
charmap [5551:5544]  = 8'b00010000;
charmap [5559:5552]  = 8'b00010000;
charmap [5567:5560]  = 8'b00000000;
charmap [5575:5568]  = 8'b10000010;
charmap [5583:5576]  = 8'b10000010;
charmap [5591:5584]  = 8'b10000010;
charmap [5599:5592]  = 8'b01010100;
charmap [5607:5600]  = 8'b01010100;
charmap [5615:5608]  = 8'b00101000;
charmap [5623:5616]  = 8'b00101000;
charmap [5631:5624]  = 8'b00000000;
charmap [5639:5632]  = 8'b01000100;
charmap [5647:5640]  = 8'b01000100;
charmap [5655:5648]  = 8'b00101000;
charmap [5663:5656]  = 8'b00010000;
charmap [5671:5664]  = 8'b00101000;
charmap [5679:5672]  = 8'b01000100;
charmap [5687:5680]  = 8'b01000100;
charmap [5695:5688]  = 8'b00000000;
charmap [5703:5696]  = 8'b01000100;
charmap [5711:5704]  = 8'b01000100;
charmap [5719:5712]  = 8'b00101000;
charmap [5727:5720]  = 8'b00010000;
charmap [5735:5728]  = 8'b00010000;
charmap [5743:5736]  = 8'b00010000;
charmap [5751:5744]  = 8'b00010000;
charmap [5759:5752]  = 8'b00000000;
charmap [5767:5760]  = 8'b01111100;
charmap [5775:5768]  = 8'b01000000;
charmap [5783:5776]  = 8'b00100000;
charmap [5791:5784]  = 8'b00010000;
charmap [5799:5792]  = 8'b00001000;
charmap [5807:5800]  = 8'b00000100;
charmap [5815:5808]  = 8'b01111100;
charmap [5823:5816]  = 8'b00000000;
charmap [5831:5824]  = 8'b00111000;
charmap [5839:5832]  = 8'b00001000;
charmap [5847:5840]  = 8'b00001000;
charmap [5855:5848]  = 8'b00001000;
charmap [5863:5856]  = 8'b00001000;
charmap [5871:5864]  = 8'b00001000;
charmap [5879:5872]  = 8'b00111000;
charmap [5887:5880]  = 8'b00000000;
charmap [5895:5888]  = 8'b00000010;
charmap [5903:5896]  = 8'b00000100;
charmap [5911:5904]  = 8'b00001000;
charmap [5919:5912]  = 8'b00010000;
charmap [5927:5920]  = 8'b00100000;
charmap [5935:5928]  = 8'b01000000;
charmap [5943:5936]  = 8'b10000000;
charmap [5951:5944]  = 8'b00000000;
charmap [5959:5952]  = 8'b00111000;
charmap [5967:5960]  = 8'b00100000;
charmap [5975:5968]  = 8'b00100000;
charmap [5983:5976]  = 8'b00100000;
charmap [5991:5984]  = 8'b00100000;
charmap [5999:5992]  = 8'b00100000;
charmap [6007:6000]  = 8'b00111000;
charmap [6015:6008]  = 8'b00000000;
charmap [6023:6016]  = 8'b00010000;
charmap [6031:6024]  = 8'b00101000;
charmap [6039:6032]  = 8'b01000100;
charmap [6047:6040]  = 8'b00000000;
charmap [6055:6048]  = 8'b00000000;
charmap [6063:6056]  = 8'b00000000;
charmap [6071:6064]  = 8'b00000000;
charmap [6079:6072]  = 8'b00000000;
charmap [6087:6080]  = 8'b00000000;
charmap [6095:6088]  = 8'b00000000;
charmap [6103:6096]  = 8'b00000000;
charmap [6111:6104]  = 8'b00000000;
charmap [6119:6112]  = 8'b00000000;
charmap [6127:6120]  = 8'b00000000;
charmap [6135:6128]  = 8'b00000000;
charmap [6143:6136]  = 8'b11111110;
charmap [6151:6144]  = 8'b00001000;
charmap [6159:6152]  = 8'b00010000;
charmap [6167:6160]  = 8'b00000000;
charmap [6175:6168]  = 8'b00000000;
charmap [6183:6176]  = 8'b00000000;
charmap [6191:6184]  = 8'b00000000;
charmap [6199:6192]  = 8'b00000000;
charmap [6207:6200]  = 8'b00000000;
charmap [6215:6208]  = 8'b00000000;
charmap [6223:6216]  = 8'b00111000;
charmap [6231:6224]  = 8'b01000000;
charmap [6239:6232]  = 8'b01111000;
charmap [6247:6240]  = 8'b01000100;
charmap [6255:6248]  = 8'b01000100;
charmap [6263:6256]  = 8'b10111000;
charmap [6271:6264]  = 8'b00000000;
charmap [6279:6272]  = 8'b00001000;
charmap [6287:6280]  = 8'b00001000;
charmap [6295:6288]  = 8'b00111000;
charmap [6303:6296]  = 8'b01001000;
charmap [6311:6304]  = 8'b01001000;
charmap [6319:6312]  = 8'b01001000;
charmap [6327:6320]  = 8'b00110100;
charmap [6335:6328]  = 8'b00000000;
charmap [6343:6336]  = 8'b00000000;
charmap [6351:6344]  = 8'b00000000;
charmap [6359:6352]  = 8'b00111000;
charmap [6367:6360]  = 8'b00000100;
charmap [6375:6368]  = 8'b00000100;
charmap [6383:6376]  = 8'b00000100;
charmap [6391:6384]  = 8'b00111000;
charmap [6399:6392]  = 8'b00000000;
charmap [6407:6400]  = 8'b01000000;
charmap [6415:6408]  = 8'b01000000;
charmap [6423:6416]  = 8'b01110000;
charmap [6431:6424]  = 8'b01001000;
charmap [6439:6432]  = 8'b01001000;
charmap [6447:6440]  = 8'b01001000;
charmap [6455:6448]  = 8'b10110000;
charmap [6463:6456]  = 8'b00000000;
charmap [6471:6464]  = 8'b00000000;
charmap [6479:6472]  = 8'b00000000;
charmap [6487:6480]  = 8'b00111000;
charmap [6495:6488]  = 8'b01000100;
charmap [6503:6496]  = 8'b01111100;
charmap [6511:6504]  = 8'b00000100;
charmap [6519:6512]  = 8'b00111000;
charmap [6527:6520]  = 8'b00000000;
charmap [6535:6528]  = 8'b00110000;
charmap [6543:6536]  = 8'b01001000;
charmap [6551:6544]  = 8'b00001000;
charmap [6559:6552]  = 8'b00011100;
charmap [6567:6560]  = 8'b00001000;
charmap [6575:6568]  = 8'b00001000;
charmap [6583:6576]  = 8'b00001000;
charmap [6591:6584]  = 8'b00000000;
charmap [6599:6592]  = 8'b00000000;
charmap [6607:6600]  = 8'b00000000;
charmap [6615:6608]  = 8'b10111000;
charmap [6623:6616]  = 8'b01000100;
charmap [6631:6624]  = 8'b01000100;
charmap [6639:6632]  = 8'b01111000;
charmap [6647:6640]  = 8'b01000000;
charmap [6655:6648]  = 8'b00111000;
charmap [6663:6656]  = 8'b00000100;
charmap [6671:6664]  = 8'b00000100;
charmap [6679:6672]  = 8'b00110100;
charmap [6687:6680]  = 8'b01001100;
charmap [6695:6688]  = 8'b01000100;
charmap [6703:6696]  = 8'b01000100;
charmap [6711:6704]  = 8'b01000100;
charmap [6719:6712]  = 8'b00000000;
charmap [6727:6720]  = 8'b00000000;
charmap [6735:6728]  = 8'b00010000;
charmap [6743:6736]  = 8'b00000000;
charmap [6751:6744]  = 8'b00010000;
charmap [6759:6752]  = 8'b00010000;
charmap [6767:6760]  = 8'b00010000;
charmap [6775:6768]  = 8'b00010000;
charmap [6783:6776]  = 8'b00000000;
charmap [6791:6784]  = 8'b00000000;
charmap [6799:6792]  = 8'b00010000;
charmap [6807:6800]  = 8'b00000000;
charmap [6815:6808]  = 8'b00010000;
charmap [6823:6816]  = 8'b00010000;
charmap [6831:6824]  = 8'b00010000;
charmap [6839:6832]  = 8'b00010000;
charmap [6847:6840]  = 8'b00001100;
charmap [6855:6848]  = 8'b00000100;
charmap [6863:6856]  = 8'b00000100;
charmap [6871:6864]  = 8'b00100100;
charmap [6879:6872]  = 8'b00010100;
charmap [6887:6880]  = 8'b00001100;
charmap [6895:6888]  = 8'b00010100;
charmap [6903:6896]  = 8'b00100100;
charmap [6911:6904]  = 8'b00000000;
charmap [6919:6912]  = 8'b00011000;
charmap [6927:6920]  = 8'b00010000;
charmap [6935:6928]  = 8'b00010000;
charmap [6943:6936]  = 8'b00010000;
charmap [6951:6944]  = 8'b00010000;
charmap [6959:6952]  = 8'b00010000;
charmap [6967:6960]  = 8'b00010000;
charmap [6975:6968]  = 8'b00000000;
charmap [6983:6976]  = 8'b00000000;
charmap [6991:6984]  = 8'b00000000;
charmap [6999:6992]  = 8'b01101101;
charmap [7007:7000]  = 8'b10010010;
charmap [7015:7008]  = 8'b10010010;
charmap [7023:7016]  = 8'b10000010;
charmap [7031:7024]  = 8'b10000010;
charmap [7039:7032]  = 8'b00000000;
charmap [7047:7040]  = 8'b00000000;
charmap [7055:7048]  = 8'b00000000;
charmap [7063:7056]  = 8'b00110100;
charmap [7071:7064]  = 8'b01001000;
charmap [7079:7072]  = 8'b01001000;
charmap [7087:7080]  = 8'b01001000;
charmap [7095:7088]  = 8'b01001000;
charmap [7103:7096]  = 8'b00000000;
charmap [7111:7104]  = 8'b00000000;
charmap [7119:7112]  = 8'b00000000;
charmap [7127:7120]  = 8'b00111000;
charmap [7135:7128]  = 8'b01000100;
charmap [7143:7136]  = 8'b01000100;
charmap [7151:7144]  = 8'b01000100;
charmap [7159:7152]  = 8'b00111000;
charmap [7167:7160]  = 8'b00000000;
charmap [7175:7168]  = 8'b00000000;
charmap [7183:7176]  = 8'b00000000;
charmap [7191:7184]  = 8'b00110100;
charmap [7199:7192]  = 8'b01001000;
charmap [7207:7200]  = 8'b01001000;
charmap [7215:7208]  = 8'b00111000;
charmap [7223:7216]  = 8'b00001000;
charmap [7231:7224]  = 8'b00001000;
charmap [7239:7232]  = 8'b00000000;
charmap [7247:7240]  = 8'b00000000;
charmap [7255:7248]  = 8'b01011000;
charmap [7263:7256]  = 8'b00100100;
charmap [7271:7264]  = 8'b00100100;
charmap [7279:7272]  = 8'b00111000;
charmap [7287:7280]  = 8'b00100000;
charmap [7295:7288]  = 8'b00100000;
charmap [7303:7296]  = 8'b00000000;
charmap [7311:7304]  = 8'b00000000;
charmap [7319:7312]  = 8'b00110100;
charmap [7327:7320]  = 8'b00001100;
charmap [7335:7328]  = 8'b00000100;
charmap [7343:7336]  = 8'b00000100;
charmap [7351:7344]  = 8'b00000100;
charmap [7359:7352]  = 8'b00000000;
charmap [7367:7360]  = 8'b00000000;
charmap [7375:7368]  = 8'b00000000;
charmap [7383:7376]  = 8'b00111000;
charmap [7391:7384]  = 8'b00000100;
charmap [7399:7392]  = 8'b00011000;
charmap [7407:7400]  = 8'b00100000;
charmap [7415:7408]  = 8'b00011100;
charmap [7423:7416]  = 8'b00000000;
charmap [7431:7424]  = 8'b00000000;
charmap [7439:7432]  = 8'b00010000;
charmap [7447:7440]  = 8'b00111000;
charmap [7455:7448]  = 8'b00010000;
charmap [7463:7456]  = 8'b00010000;
charmap [7471:7464]  = 8'b00010000;
charmap [7479:7472]  = 8'b00010000;
charmap [7487:7480]  = 8'b00000000;
charmap [7495:7488]  = 8'b00000000;
charmap [7503:7496]  = 8'b00000000;
charmap [7511:7504]  = 8'b00100100;
charmap [7519:7512]  = 8'b00100100;
charmap [7527:7520]  = 8'b00100100;
charmap [7535:7528]  = 8'b00100100;
charmap [7543:7536]  = 8'b01011000;
charmap [7551:7544]  = 8'b00000000;
charmap [7559:7552]  = 8'b00000000;
charmap [7567:7560]  = 8'b00000000;
charmap [7575:7568]  = 8'b01000100;
charmap [7583:7576]  = 8'b01000100;
charmap [7591:7584]  = 8'b01000100;
charmap [7599:7592]  = 8'b00101000;
charmap [7607:7600]  = 8'b00010000;
charmap [7615:7608]  = 8'b00000000;
charmap [7623:7616]  = 8'b00000000;
charmap [7631:7624]  = 8'b00000000;
charmap [7639:7632]  = 8'b10000010;
charmap [7647:7640]  = 8'b10000010;
charmap [7655:7648]  = 8'b10010010;
charmap [7663:7656]  = 8'b10101010;
charmap [7671:7664]  = 8'b01000100;
charmap [7679:7672]  = 8'b00000000;
charmap [7687:7680]  = 8'b00000000;
charmap [7695:7688]  = 8'b00000000;
charmap [7703:7696]  = 8'b01000100;
charmap [7711:7704]  = 8'b00101000;
charmap [7719:7712]  = 8'b00010000;
charmap [7727:7720]  = 8'b00101000;
charmap [7735:7728]  = 8'b01000100;
charmap [7743:7736]  = 8'b00000000;
charmap [7751:7744]  = 8'b00000000;
charmap [7759:7752]  = 8'b00000000;
charmap [7767:7760]  = 8'b01001000;
charmap [7775:7768]  = 8'b01001000;
charmap [7783:7776]  = 8'b01001000;
charmap [7791:7784]  = 8'b01110000;
charmap [7799:7792]  = 8'b01000000;
charmap [7807:7800]  = 8'b00111000;
charmap [7815:7808]  = 8'b00000000;
charmap [7823:7816]  = 8'b00000000;
charmap [7831:7824]  = 8'b00111100;
charmap [7839:7832]  = 8'b00100000;
charmap [7847:7840]  = 8'b00010000;
charmap [7855:7848]  = 8'b00001000;
charmap [7863:7856]  = 8'b00111100;
charmap [7871:7864]  = 8'b00000000;
charmap [7879:7872]  = 8'b00110000;
charmap [7887:7880]  = 8'b00001000;
charmap [7895:7888]  = 8'b00001000;
charmap [7903:7896]  = 8'b00000100;
charmap [7911:7904]  = 8'b00001000;
charmap [7919:7912]  = 8'b00001000;
charmap [7927:7920]  = 8'b00110000;
charmap [7935:7928]  = 8'b00000000;
charmap [7943:7936]  = 8'b00010000;
charmap [7951:7944]  = 8'b00010000;
charmap [7959:7952]  = 8'b00010000;
charmap [7967:7960]  = 8'b00010000;
charmap [7975:7968]  = 8'b00010000;
charmap [7983:7976]  = 8'b00010000;
charmap [7991:7984]  = 8'b00010000;
charmap [7999:7992]  = 8'b00000000;
charmap [8007:8000]  = 8'b00001100;
charmap [8015:8008]  = 8'b00010000;
charmap [8023:8016]  = 8'b00010000;
charmap [8031:8024]  = 8'b00100000;
charmap [8039:8032]  = 8'b00010000;
charmap [8047:8040]  = 8'b00010000;
charmap [8055:8048]  = 8'b00001100;
charmap [8063:8056]  = 8'b00000000;
charmap [8071:8064]  = 8'b00000000;
charmap [8079:8072]  = 8'b00000000;
charmap [8087:8080]  = 8'b00001100;
charmap [8095:8088]  = 8'b10010010;
charmap [8103:8096]  = 8'b01100000;
charmap [8111:8104]  = 8'b00000000;
charmap [8119:8112]  = 8'b00000000;
charmap [8127:8120]  = 8'b00000000;
charmap [8135:8128]  = 8'b00000000;
charmap [8143:8136]  = 8'b00000000;
charmap [8151:8144]  = 8'b00000000;
charmap [8159:8152]  = 8'b00000000;
charmap [8167:8160]  = 8'b00000000;
charmap [8175:8168]  = 8'b00000000;
charmap [8183:8176]  = 8'b00000000;
charmap [8191:8184]  = 8'b00000000;

end


always @( posedge CLK_108MHz or posedge reset)
begin
	if(reset)
	begin
		hsync_out <= 1'b0;
		vsync_out <= 1'b0;
		de_out 		<= 1'b0;
		color_out <= 8'h00;
	end
	else
	begin
		hsync_out <= hsync_in;
		vsync_out <= vsync_in;
		de_out 		<= de_in;
		color_out <= color_in;
	end
end
	


// look up the pixel value

always @ (posedge CLK_108MHz)
begin
	if(reset)
	begin
		pixel_out <= pixel_out;
	end
	else
	begin
		pixel_out <= de_in ? charmap[ {character_in, vctr_in, hctr_in} ] : 1'b0;
	end
end

endmodule
